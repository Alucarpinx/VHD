LIBRARY IEEE;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;            
USE ieee.std_logic_unsigned.all;

ENTITY 




Component mux is 
	      ( )
			
END Component; 

Component delay_unit is 
	      ( )
			
END Component; 

Component shifter is 
	      ( )
			
END Component; 